/*
 This module is testbench for or1200_ctrl.v
 or1200_ctrl.v is modified for keccak.

 */

//`timescale 1ns / 1ps
`define P 200



module test_sign;

   // Inputs
   reg clk;
   reg rst;
   reg [511:0] message;
   // Outputs
   wire [232:0] sign_u;
   wire [232:0] sign_v;
   wire done;
   // Instantiate the Unit Under Test (UUT)
   ecdsa_sign ed1(
    .clk(clk),
    .nrst(rst),
    .message(message),
    .sign_u(sign_u),
    .sign_v(sign_v),
    .done(done)
      );
   initial begin
      // Initialize Inputs
      clk = 0;
      rst = 0;
message = 512'b01100001_01100010_01100011_01100100_01100010_01100011_01100100_01100101_01100011_01100100_01100101_01100110_01100100_01100101_01100110_01100111_01100101_01100110_01100111_01101000_01100110_01100111_01101000_01101001_01100111_01101000_01101001_01101010_01101000_01101001_01101010_01101011_01101001_01101010_01101011_01101100_01101010_01101011_01101100_01101101_01101011_01101100_01101101_01101110_01101100_01101101_01101110_01101111_01101101_01101110_01101111_01110000_01101110_01101111_01110000_01110001_01110001_01110001_01110001_01110001_01110001_01110001_01110001_01110001;

      // Wait 100 ns for global reset to finish
      #100;

      // Add stimulus here
      @ (negedge clk);

      //test vector
  		#10	rst = 1'b0;
		#110 	rst = 1'b1;
		#3080 rst = 1'b0;
		#100 rst = 1'b1;
		#3000 rst = 1'b0;
      //message = 512'h FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF;
      #(`P);
      //message = 512'h 000a02b784e94a02b733e94a02baa4e33a02b784e33a02b784e94a02444;
      #100 message = 512'b01100001_01100010_01100011_01100100_01100010_01100011_01100100_01100101_01100011_01100100_01100101_01100110_01100100_01100101_01100110_01100111_01100101_01100110_01100111_01101000_01100110_01100111_01101000_01101001_01100111_01101000_01101001_01101010_01101000_01101001_01101010_01101011_01101001_01101010_01101011_01101100_01101010_01101011_01101100_01101101_01101011_01101100_01101101_01101110_01101100_01101101_01101110_01101111_01101101_01101110_01101111_01110000_01101110_01101111_01110000_01110001_01110001_01110001_01110001_01110001_01110001_01110001_01110001_01110001;
    #200 rst = 1'b1;
    #10000000 rst = 1'b0;
       end
   //always #(`P/2) clk = ~ clk;
always #100 clk = ~ clk;

   task error;
      begin
         $display("E");
         $finish;
      end
   endtask


endmodule

`undef P
